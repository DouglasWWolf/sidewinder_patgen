
//================================================================================================
//    Date         Version     Who  Changes
// -----------------------------------------------------------------------------------------------
// 25-Oct-2023     1.0.1       DWW  Initial creation
//
// 06-Dec-2023     1.0.2       DWW  Fixed bug loading FIFO #2, added signal added "new_job"
//================================================================================================
localparam VERSION_MAJOR = 1;
localparam VERSION_MINOR = 0;
localparam VERSION_BUILD = 2;
localparam VERSION_RCAND = 0;

localparam VERSION_DAY   = 06;
localparam VERSION_MONTH = 12;
localparam VERSION_YEAR  = 2023;
